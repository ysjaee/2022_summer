module ripp