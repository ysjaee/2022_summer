module binary_counter()