module Twos_Complement_Substraction()
