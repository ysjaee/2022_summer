module testbench();
    reg [31:0]x;
    reg [31:0]y;
    reg ci;
    wire co;
    wire [31:0]res;


    Ripple_carry_addition Rcat(.x(x),.y(y),.ci(ci),.co(co),.res(res));

    initial begin
        x = 32'h00000000; y = 32'h00000000; ci = 1'b0;
        #3 x = 32'h00000001; y = 32'h00000001; ci = 1'b1;
        #6 x = 32'h00000010; y = 32'h00000010; ci = 1'b1;
        #9 x = 32'h00000010; y = 32'h00000010; ci = 1'b0;
        #12 x = 32'h00000011; y = 32'h00000011; ci = 1'b1;
        #15 x = 32'h00000011; y = 32'h00000011; ci = 1'b0;        
        #21 x = 32'h00000011; y = 32'h00000011; ci = 1'b0;
        #24 x = 32'h00000100; y = 32'h00000100; ci = 1'b1;
        #27 x = 32'h00000100; y = 32'h00000100; ci = 1'b0;
        #30 x = 32'h00001000; y = 32'h00001000; ci = 1'b1;
        #33 x = 32'h00001000; y = 32'h00001000; ci = 1'b0;
        #36 x = 32'h10001000; y = 32'h10001000; ci = 1'b1;
        #60 $stop;
    end
endmodule